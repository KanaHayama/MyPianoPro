library verilog;
use verilog.vl_types.all;
entity ToneGenerator_vlg_vec_tst is
end ToneGenerator_vlg_vec_tst;
