library verilog;
use verilog.vl_types.all;
entity FreqChange_vlg_vec_tst is
end FreqChange_vlg_vec_tst;
